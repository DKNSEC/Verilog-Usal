module prueba;

integer a;  
integer b;

initial

	begin

	a = 1;
	b = 'b1001;

	/*--------------------------------------------------------------------------------*/

	$display("%d", a);
	$display("%d", b);

	end

endmodule