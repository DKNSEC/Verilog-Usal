/* Programa de ejemplo: hello.v */

module hello;

  initial

    $display("Hola, mundo\nHola, mundo \n");

endmodule