module prueba;

initial
	begin

	$display("Estamos recordando como programar con Verilog");

	end
endmodule