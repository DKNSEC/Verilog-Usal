/* Programa de ejemplo: hello.v */

module hello;

  initial
    // Imprimimos el mensaje y un salto de lInea
    $display("Hola, mundo\n");

endmodule
